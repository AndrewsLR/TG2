A equação é :((a+b)*(c+d))
M1 n1 a GND GND nfet
M2 GND b n1 GND nfet
M3 n2 c n1 GND nfet
M4 n1 d n2 GND nfet
M5 VDD a n3 VDD pfet
M6 n3 b n2 VDD pfet
M7 VDD c n5 VDD pfet
M8 n5 d n2 VDD pfet
M1 n1 a GND GND nfet
M2 GND b n1 GND nfet
M3 n2 c n1 GND nfet
M4 n1 d n2 GND nfet
M5 VDD a n3 VDD pfet
M6 n3 b n2 VDD pfet
M7 n5 c VDD VDD pfet
M8 n2 d n5 VDD pfet
A equação é :((a+b)*(c+d))
M1 n1 a GND GND nfet
M2 GND b n1 GND nfet
M3 n2 c n1 GND nfet
M4 n1 d n2 GND nfet
M5 VDD a n3 VDD pfet
M6 n3 b n2 VDD pfet
M7 VDD c n5 VDD pfet
M8 n5 d n2 VDD pfet
M1 n1 a GND GND nfet
M2 GND b n1 GND nfet
M3 n2 c n1 GND nfet
M4 n1 d n2 GND nfet
M5 VDD a n3 VDD pfet
M6 n3 b n2 VDD pfet
M7 n5 c VDD VDD pfet
M8 n2 d n5 VDD pfet
