A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :CONST0
A equação é :CONST1
A equação é :a
A equação é :(a*b)
M1 n1 a GND GND nfet
M2 n2 b n1 GND nfet
M3 n2 a VDD VDD pfet
M4 n2 b VDD VDD pfet
A equação é :(a*(b+c))
M1 n1 b GND GND nfet
M2 n1 c GND GND nfet
M3 n2 a n1 GND nfet
M4 n3 b VDD VDD pfet
M5 n2 c n3 VDD pfet
M6 n2 a VDD VDD pfet
A equação é :(a*(b+c*d))
M1 n1 c GND GND nfet
M2 n2 d n1 GND nfet
M3 n2 b GND GND nfet
M4 n3 a n2 GND nfet
M5 n4 c VDD VDD pfet
M6 n4 d VDD VDD pfet
M7 n3 b n4 VDD pfet
M8 n3 a VDD VDD pfet
A equação é :(a*(b+c*(d+e)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n2 c n1 GND nfet
M4 n2 b GND GND nfet
M5 n3 a n2 GND nfet
M6 n4 d VDD VDD pfet
M7 n5 e n4 VDD pfet
M8 n5 c VDD VDD pfet
M9 n3 b n5 VDD pfet
M10 n3 a VDD VDD pfet
A equação é :(a*(b+c*(d+e*f)))
M1 n1 e GND GND nfet
M2 n2 f n1 GND nfet
M3 n2 d GND GND nfet
M4 n3 c n2 GND nfet
M5 n3 b GND GND nfet
M6 n4 a n3 GND nfet
M7 n5 e VDD VDD pfet
M8 n5 f VDD VDD pfet
M9 n6 d n5 VDD pfet
M10 n6 c VDD VDD pfet
M11 n4 b n6 VDD pfet
M12 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+e*(f+g))))
M1 n1 f GND GND nfet
M2 n1 g GND GND nfet
M3 n2 e n1 GND nfet
M4 n2 d GND GND nfet
M5 n3 c n2 GND nfet
M6 n3 b GND GND nfet
M7 n4 a n3 GND nfet
M8 n5 f VDD VDD pfet
M9 n6 g n5 VDD pfet
M10 n6 e VDD VDD pfet
M11 n7 d n6 VDD pfet
M12 n7 c VDD VDD pfet
M13 n4 b n7 VDD pfet
M14 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+(e+f)*(g+h))))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n3 c n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 e VDD VDD pfet
M10 n4 f n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 h n7 VDD pfet
M13 n9 d n4 VDD pfet
M14 n9 c VDD VDD pfet
M15 n4 b n9 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d*e+f*g)))
M1 n1 d GND GND nfet
M2 n6 e n1 GND nfet
M3 n3 f GND GND nfet
M4 n6 g n3 GND nfet
M5 n5 c n6 GND nfet
M6 n5 b GND GND nfet
M7 n6 a n5 GND nfet
M8 n7 d VDD VDD pfet
M9 n7 e VDD VDD pfet
M10 n8 f n7 VDD pfet
M11 n8 g n7 VDD pfet
M12 n8 c VDD VDD pfet
M13 n6 b n8 VDD pfet
M14 n6 a VDD VDD pfet
A equação é :(a*(b+c*(d*e+f*(g+h))))
M1 n1 d GND GND nfet
M2 n6 e n1 GND nfet
M3 n3 g GND GND nfet
M4 n3 h GND GND nfet
M5 n6 f n3 GND nfet
M6 n5 c n6 GND nfet
M7 n5 b GND GND nfet
M8 n6 a n5 GND nfet
M9 n7 d VDD VDD pfet
M10 n7 e VDD VDD pfet
M11 n8 g n7 VDD pfet
M12 n9 h n8 VDD pfet
M13 n9 f n7 VDD pfet
M14 n9 c VDD VDD pfet
M15 n6 b n9 VDD pfet
M16 n6 a VDD VDD pfet
A equação é :(a*(b+c*(d*e+(f+g)*(h+i))))
M1 n1 f GND GND nfet
M2 n1 g GND GND nfet
M3 n6 h n1 GND nfet
M4 n6 i n1 GND nfet
M5 n3 d GND GND nfet
M6 n6 e n3 GND nfet
M7 n5 c n6 GND nfet
M8 n5 b GND GND nfet
M9 n6 a n5 GND nfet
M10 n7 f VDD VDD pfet
M11 n6 g n7 VDD pfet
M12 n9 h VDD VDD pfet
M13 n6 i n9 VDD pfet
M14 n11 d n6 VDD pfet
M15 n11 e n6 VDD pfet
M16 n11 c VDD VDD pfet
M17 n6 b n11 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b+c*(d+e+f)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n1 f GND GND nfet
M4 n2 c n1 GND nfet
M5 n2 b GND GND nfet
M6 n3 a n2 GND nfet
M7 n4 d VDD VDD pfet
M8 n5 e n4 VDD pfet
M9 n6 f n5 VDD pfet
M10 n6 c VDD VDD pfet
M11 n3 b n6 VDD pfet
M12 n3 a VDD VDD pfet
A equação é :(a*(b+c*(d+e+f*g)))
M1 n5 d GND GND nfet
M2 n5 e GND GND nfet
M3 n2 f GND GND nfet
M4 n5 g n2 GND nfet
M5 n4 c n5 GND nfet
M6 n4 b GND GND nfet
M7 n5 a n4 GND nfet
M8 n6 d VDD VDD pfet
M9 n7 e n6 VDD pfet
M10 n8 f n7 VDD pfet
M11 n8 g n7 VDD pfet
M12 n8 c VDD VDD pfet
M13 n5 b n8 VDD pfet
M14 n5 a VDD VDD pfet
A equação é :(a*(b+c*(d+e*f+g*h)))
M1 n1 e GND GND nfet
M2 n6 f n1 GND nfet
M3 n6 d GND GND nfet
M4 n3 g GND GND nfet
M5 n6 h n3 GND nfet
M6 n5 c n6 GND nfet
M7 n5 b GND GND nfet
M8 n6 a n5 GND nfet
M9 n7 e VDD VDD pfet
M10 n7 f VDD VDD pfet
M11 n8 d n7 VDD pfet
M12 n9 g n8 VDD pfet
M13 n9 h n8 VDD pfet
M14 n9 c VDD VDD pfet
M15 n6 b n9 VDD pfet
M16 n6 a VDD VDD pfet
A equação é :(a*(b+c*(d*e+f*g+h*i)))
M1 n1 d GND GND nfet
M2 n8 e n1 GND nfet
M3 n3 f GND GND nfet
M4 n8 g n3 GND nfet
M5 n5 h GND GND nfet
M6 n8 i n5 GND nfet
M7 n7 c n8 GND nfet
M8 n7 b GND GND nfet
M9 n8 a n7 GND nfet
M10 n9 d VDD VDD pfet
M11 n9 e VDD VDD pfet
M12 n10 f n9 VDD pfet
M13 n10 g n9 VDD pfet
M14 n11 h n10 VDD pfet
M15 n11 i n10 VDD pfet
M16 n11 c VDD VDD pfet
M17 n8 b n11 VDD pfet
M18 n8 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+f)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 e n1 GND nfet
M4 n2 f n1 GND nfet
M5 n2 b GND GND nfet
M6 n3 a n2 GND nfet
M7 n4 c VDD VDD pfet
M8 n3 d n4 VDD pfet
M9 n6 e VDD VDD pfet
M10 n3 f n6 VDD pfet
M11 n3 b n3 VDD pfet
M12 n3 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+f*g)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 f n1 GND nfet
M4 n3 g n2 GND nfet
M5 n3 e n1 GND nfet
M6 n3 b GND GND nfet
M7 n4 a n3 GND nfet
M8 n5 c VDD VDD pfet
M9 n4 d n5 VDD pfet
M10 n7 f VDD VDD pfet
M11 n7 g VDD VDD pfet
M12 n4 e n7 VDD pfet
M13 n4 b n4 VDD pfet
M14 n4 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+f*(g+h))))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n3 f n2 GND nfet
M6 n3 e n1 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 c VDD VDD pfet
M10 n4 d n5 VDD pfet
M11 n7 g VDD VDD pfet
M12 n8 h n7 VDD pfet
M13 n8 f VDD VDD pfet
M14 n4 e n8 VDD pfet
M15 n4 b n4 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+(f+g)*(h+i))))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 f n1 GND nfet
M4 n2 g n1 GND nfet
M5 n3 h n2 GND nfet
M6 n3 i n2 GND nfet
M7 n3 e n1 GND nfet
M8 n3 b GND GND nfet
M9 n4 a n3 GND nfet
M10 n5 c VDD VDD pfet
M11 n4 d n5 VDD pfet
M12 n7 f VDD VDD pfet
M13 n4 g n7 VDD pfet
M14 n9 h VDD VDD pfet
M15 n4 i n9 VDD pfet
M16 n4 e n4 VDD pfet
M17 n4 b n4 VDD pfet
M18 n4 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e*f+g*h)))
M1 n1 e GND GND nfet
M2 n6 f n1 GND nfet
M3 n3 g GND GND nfet
M4 n6 h n3 GND nfet
M5 n5 c n6 GND nfet
M6 n5 d n6 GND nfet
M7 n5 b GND GND nfet
M8 n6 a n5 GND nfet
M9 n7 e VDD VDD pfet
M10 n7 f VDD VDD pfet
M11 n6 g n7 VDD pfet
M12 n6 h n7 VDD pfet
M13 n9 c VDD VDD pfet
M14 n6 d n9 VDD pfet
M15 n6 b n6 VDD pfet
M16 n6 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e*f+g*(h+i))))
M1 n1 e GND GND nfet
M2 n6 f n1 GND nfet
M3 n3 h GND GND nfet
M4 n3 i GND GND nfet
M5 n6 g n3 GND nfet
M6 n5 c n6 GND nfet
M7 n5 d n6 GND nfet
M8 n5 b GND GND nfet
M9 n6 a n5 GND nfet
M10 n7 e VDD VDD pfet
M11 n7 f VDD VDD pfet
M12 n8 h n7 VDD pfet
M13 n6 i n8 VDD pfet
M14 n6 g n7 VDD pfet
M15 n10 c VDD VDD pfet
M16 n6 d n10 VDD pfet
M17 n6 b n6 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e*f+(g+h)*(i+j))))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n6 i n2 GND nfet
M6 n6 j n2 GND nfet
M7 n4 e n1 GND nfet
M8 n6 f n4 GND nfet
M9 n6 b GND GND nfet
M10 n6 a n6 GND nfet
M11 n7 c VDD VDD pfet
M12 n6 d n7 VDD pfet
M13 n9 g VDD VDD pfet
M14 n6 h n9 VDD pfet
M15 n11 i VDD VDD pfet
M16 n6 j n11 VDD pfet
M17 n6 e n6 VDD pfet
M18 n6 f n6 VDD pfet
M19 n6 b n6 VDD pfet
M20 n6 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+f+g)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 e n1 GND nfet
M4 n2 f n1 GND nfet
M5 n2 g n1 GND nfet
M6 n2 b GND GND nfet
M7 n3 a n2 GND nfet
M8 n4 c VDD VDD pfet
M9 n3 d n4 VDD pfet
M10 n6 e VDD VDD pfet
M11 n7 f n6 VDD pfet
M12 n3 g n7 VDD pfet
M13 n3 b n3 VDD pfet
M14 n3 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+f+g*h)))
M1 n5 e GND GND nfet
M2 n5 f GND GND nfet
M3 n2 g GND GND nfet
M4 n5 h n2 GND nfet
M5 n4 c n5 GND nfet
M6 n4 d n5 GND nfet
M7 n4 b GND GND nfet
M8 n5 a n4 GND nfet
M9 n6 e VDD VDD pfet
M10 n7 f n6 VDD pfet
M11 n5 g n7 VDD pfet
M12 n5 h n7 VDD pfet
M13 n9 c VDD VDD pfet
M14 n5 d n9 VDD pfet
M15 n5 b n5 VDD pfet
M16 n5 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+f*g+h*i)))
M1 n1 f GND GND nfet
M2 n6 g n1 GND nfet
M3 n6 e GND GND nfet
M4 n3 h GND GND nfet
M5 n6 i n3 GND nfet
M6 n5 c n6 GND nfet
M7 n5 d n6 GND nfet
M8 n5 b GND GND nfet
M9 n6 a n5 GND nfet
M10 n7 f VDD VDD pfet
M11 n7 g VDD VDD pfet
M12 n8 e n7 VDD pfet
M13 n6 h n8 VDD pfet
M14 n6 i n8 VDD pfet
M15 n10 c VDD VDD pfet
M16 n6 d n10 VDD pfet
M17 n6 b n6 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e*f+g*h+i*j)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 e n1 GND nfet
M4 n8 f n2 GND nfet
M5 n4 g n1 GND nfet
M6 n8 h n4 GND nfet
M7 n6 i n1 GND nfet
M8 n8 j n6 GND nfet
M9 n8 b GND GND nfet
M10 n8 a n8 GND nfet
M11 n9 c VDD VDD pfet
M12 n8 d n9 VDD pfet
M13 n11 e VDD VDD pfet
M14 n11 f VDD VDD pfet
M15 n12 g n11 VDD pfet
M16 n12 h n11 VDD pfet
M17 n8 i n12 VDD pfet
M18 n8 j n12 VDD pfet
M19 n8 b n8 VDD pfet
M20 n8 a VDD VDD pfet
A equação é :(a*(b+(c+d*e)*(f+g+h)))
M1 n1 d GND GND nfet
M2 n2 e n1 GND nfet
M3 n2 c GND GND nfet
M4 n3 f n2 GND nfet
M5 n3 g n2 GND nfet
M6 n3 h n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 d VDD VDD pfet
M10 n5 e VDD VDD pfet
M11 n4 c n5 VDD pfet
M12 n7 f VDD VDD pfet
M13 n8 g n7 VDD pfet
M14 n4 h n8 VDD pfet
M15 n4 b n4 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+(c+d*(e+f))*(g+h+i)))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 d n1 GND nfet
M4 n2 c GND GND nfet
M5 n3 g n2 GND nfet
M6 n3 h n2 GND nfet
M7 n3 i n2 GND nfet
M8 n3 b GND GND nfet
M9 n4 a n3 GND nfet
M10 n5 e VDD VDD pfet
M11 n6 f n5 VDD pfet
M12 n6 d VDD VDD pfet
M13 n4 c n6 VDD pfet
M14 n8 g VDD VDD pfet
M15 n9 h n8 VDD pfet
M16 n4 i n9 VDD pfet
M17 n4 b n4 VDD pfet
M18 n4 a VDD VDD pfet
A equação é :(a*(b+(c+(d+e)*(f+g))*(h+i+j)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n2 f n1 GND nfet
M4 n2 g n1 GND nfet
M5 n2 c GND GND nfet
M6 n3 h n2 GND nfet
M7 n3 i n2 GND nfet
M8 n3 j n2 GND nfet
M9 n3 b GND GND nfet
M10 n4 a n3 GND nfet
M11 n5 d VDD VDD pfet
M12 n4 e n5 VDD pfet
M13 n7 f VDD VDD pfet
M14 n4 g n7 VDD pfet
M15 n4 c n4 VDD pfet
M16 n10 h VDD VDD pfet
M17 n11 i n10 VDD pfet
M18 n4 j n11 VDD pfet
M19 n4 b n4 VDD pfet
M20 n4 a VDD VDD pfet
A equação é :(a*(b+(c*d+e*f)*(g+h+i)))
M1 n1 c GND GND nfet
M2 n6 d n1 GND nfet
M3 n3 e GND GND nfet
M4 n6 f n3 GND nfet
M5 n5 g n6 GND nfet
M6 n5 h n6 GND nfet
M7 n5 i n6 GND nfet
M8 n5 b GND GND nfet
M9 n6 a n5 GND nfet
M10 n7 c VDD VDD pfet
M11 n7 d VDD VDD pfet
M12 n6 e n7 VDD pfet
M13 n6 f n7 VDD pfet
M14 n9 g VDD VDD pfet
M15 n10 h n9 VDD pfet
M16 n6 i n10 VDD pfet
M17 n6 b n6 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b+(c*d+e*(f+g))*(h+i+j)))
M1 n1 c GND GND nfet
M2 n6 d n1 GND nfet
M3 n3 f GND GND nfet
M4 n3 g GND GND nfet
M5 n6 e n3 GND nfet
M6 n5 h n6 GND nfet
M7 n5 i n6 GND nfet
M8 n5 j n6 GND nfet
M9 n5 b GND GND nfet
M10 n6 a n5 GND nfet
M11 n7 c VDD VDD pfet
M12 n7 d VDD VDD pfet
M13 n8 f n7 VDD pfet
M14 n6 g n8 VDD pfet
M15 n6 e n7 VDD pfet
M16 n10 h VDD VDD pfet
M17 n11 i n10 VDD pfet
M18 n6 j n11 VDD pfet
M19 n6 b n6 VDD pfet
M20 n6 a VDD VDD pfet
A equação é :(a*(b+(c*d+(e+f)*(g+h))*(i+j+k)))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n6 g n1 GND nfet
M4 n6 h n1 GND nfet
M5 n3 c GND GND nfet
M6 n6 d n3 GND nfet
M7 n5 i n6 GND nfet
M8 n5 j n6 GND nfet
M9 n5 k n6 GND nfet
M10 n5 b GND GND nfet
M11 n6 a n5 GND nfet
M12 n7 e VDD VDD pfet
M13 n6 f n7 VDD pfet
M14 n9 g VDD VDD pfet
M15 n6 h n9 VDD pfet
M16 n6 c n6 VDD pfet
M17 n6 d n6 VDD pfet
M18 n12 i VDD VDD pfet
M19 n13 j n12 VDD pfet
M20 n6 k n13 VDD pfet
M21 n6 b n6 VDD pfet
M22 n6 a VDD VDD pfet
A equação é :(a*(b+(c+d+e)*(f+g+h)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n1 e GND GND nfet
M4 n2 f n1 GND nfet
M5 n2 g n1 GND nfet
M6 n2 h n1 GND nfet
M7 n2 b GND GND nfet
M8 n3 a n2 GND nfet
M9 n4 c VDD VDD pfet
M10 n5 d n4 VDD pfet
M11 n3 e n5 VDD pfet
M12 n7 f VDD VDD pfet
M13 n8 g n7 VDD pfet
M14 n3 h n8 VDD pfet
M15 n3 b n3 VDD pfet
M16 n3 a VDD VDD pfet
A equação é :(a*(b+(c+d+e)*(f+g+h*i)))
M1 n5 f GND GND nfet
M2 n5 g GND GND nfet
M3 n2 h GND GND nfet
M4 n5 i n2 GND nfet
M5 n4 c n5 GND nfet
M6 n4 d n5 GND nfet
M7 n4 e n5 GND nfet
M8 n4 b GND GND nfet
M9 n5 a n4 GND nfet
M10 n6 f VDD VDD pfet
M11 n7 g n6 VDD pfet
M12 n5 h n7 VDD pfet
M13 n5 i n7 VDD pfet
M14 n9 c VDD VDD pfet
M15 n10 d n9 VDD pfet
M16 n5 e n10 VDD pfet
M17 n5 b n5 VDD pfet
M18 n5 a VDD VDD pfet
A equação é :(a*(b+(c+d+e)*(f+g*h+i*j)))
M1 n1 g GND GND nfet
M2 n6 h n1 GND nfet
M3 n6 f GND GND nfet
M4 n3 i GND GND nfet
M5 n6 j n3 GND nfet
M6 n5 c n6 GND nfet
M7 n5 d n6 GND nfet
M8 n5 e n6 GND nfet
M9 n5 b GND GND nfet
M10 n6 a n5 GND nfet
M11 n7 g VDD VDD pfet
M12 n7 h VDD VDD pfet
M13 n8 f n7 VDD pfet
M14 n6 i n8 VDD pfet
M15 n6 j n8 VDD pfet
M16 n10 c VDD VDD pfet
M17 n11 d n10 VDD pfet
M18 n6 e n11 VDD pfet
M19 n6 b n6 VDD pfet
M20 n6 a VDD VDD pfet
A equação é :(a*(b+(c+d+e)*(f*g+h*i+j*k)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n1 e GND GND nfet
M4 n2 f n1 GND nfet
M5 n8 g n2 GND nfet
M6 n4 h n1 GND nfet
M7 n8 i n4 GND nfet
M8 n6 j n1 GND nfet
M9 n8 k n6 GND nfet
M10 n8 b GND GND nfet
M11 n8 a n8 GND nfet
M12 n9 c VDD VDD pfet
M13 n10 d n9 VDD pfet
M14 n8 e n10 VDD pfet
M15 n12 f VDD VDD pfet
M16 n12 g VDD VDD pfet
M17 n13 h n12 VDD pfet
M18 n13 i n12 VDD pfet
M19 n8 j n13 VDD pfet
M20 n8 k n13 VDD pfet
M21 n8 b n8 VDD pfet
M22 n8 a VDD VDD pfet
A equação é :(a*(b+c*d*e))
M1 n1 c GND GND nfet
M2 n2 d n1 GND nfet
M3 n3 e n2 GND nfet
M4 n3 b GND GND nfet
M5 n4 a n3 GND nfet
M6 n5 c VDD VDD pfet
M7 n5 d VDD VDD pfet
M8 n5 e VDD VDD pfet
M9 n4 b n5 VDD pfet
M10 n4 a VDD VDD pfet
A equação é :(a*(b+c*d*(e+f)))
M1 n1 c GND GND nfet
M2 n2 d n1 GND nfet
M3 n3 e n2 GND nfet
M4 n3 f n2 GND nfet
M5 n3 b GND GND nfet
M6 n4 a n3 GND nfet
M7 n4 c VDD VDD pfet
M8 n4 d VDD VDD pfet
M9 n6 e VDD VDD pfet
M10 n4 f n6 VDD pfet
M11 n4 b n4 VDD pfet
M12 n4 a VDD VDD pfet
A equação é :(a*(b+c*d*(e+f+g)))
M1 n1 c GND GND nfet
M2 n2 d n1 GND nfet
M3 n3 e n2 GND nfet
M4 n3 f n2 GND nfet
M5 n3 g n2 GND nfet
M6 n3 b GND GND nfet
M7 n4 a n3 GND nfet
M8 n4 c VDD VDD pfet
M9 n4 d VDD VDD pfet
M10 n6 e VDD VDD pfet
M11 n7 f n6 VDD pfet
M12 n4 g n7 VDD pfet
M13 n4 b n4 VDD pfet
M14 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+e)*(f+g)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n2 c n1 GND nfet
M4 n3 f n2 GND nfet
M5 n3 g n2 GND nfet
M6 n3 b GND GND nfet
M7 n4 a n3 GND nfet
M8 n5 d VDD VDD pfet
M9 n4 e n5 VDD pfet
M10 n4 c VDD VDD pfet
M11 n7 f VDD VDD pfet
M12 n4 g n7 VDD pfet
M13 n4 b n4 VDD pfet
M14 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+e)*(f+g+h)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n2 c n1 GND nfet
M4 n3 f n2 GND nfet
M5 n3 g n2 GND nfet
M6 n3 h n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 d VDD VDD pfet
M10 n4 e n5 VDD pfet
M11 n4 c VDD VDD pfet
M12 n7 f VDD VDD pfet
M13 n8 g n7 VDD pfet
M14 n4 h n8 VDD pfet
M15 n4 b n4 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+c*(d+e+f)*(g+h+i)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n1 f GND GND nfet
M4 n2 c n1 GND nfet
M5 n3 g n2 GND nfet
M6 n3 h n2 GND nfet
M7 n3 i n2 GND nfet
M8 n3 b GND GND nfet
M9 n4 a n3 GND nfet
M10 n5 d VDD VDD pfet
M11 n6 e n5 VDD pfet
M12 n4 f n6 VDD pfet
M13 n4 c VDD VDD pfet
M14 n8 g VDD VDD pfet
M15 n9 h n8 VDD pfet
M16 n4 i n9 VDD pfet
M17 n4 b n4 VDD pfet
M18 n4 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+f)*(g+h)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 e n1 GND nfet
M4 n2 f n1 GND nfet
M5 n3 g n2 GND nfet
M6 n3 h n2 GND nfet
M7 n3 b GND GND nfet
M8 n4 a n3 GND nfet
M9 n5 c VDD VDD pfet
M10 n4 d n5 VDD pfet
M11 n7 e VDD VDD pfet
M12 n4 f n7 VDD pfet
M13 n9 g VDD VDD pfet
M14 n4 h n9 VDD pfet
M15 n4 b n4 VDD pfet
M16 n4 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+f)*(g+h+i)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 e n1 GND nfet
M4 n2 f n1 GND nfet
M5 n3 g n2 GND nfet
M6 n3 h n2 GND nfet
M7 n3 i n2 GND nfet
M8 n3 b GND GND nfet
M9 n4 a n3 GND nfet
M10 n5 c VDD VDD pfet
M11 n4 d n5 VDD pfet
M12 n7 e VDD VDD pfet
M13 n4 f n7 VDD pfet
M14 n9 g VDD VDD pfet
M15 n10 h n9 VDD pfet
M16 n4 i n10 VDD pfet
M17 n4 b n4 VDD pfet
M18 n4 a VDD VDD pfet
A equação é :(a*(b+(c+d)*(e+f+g)*(h+i+j)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n2 e n1 GND nfet
M4 n2 f n1 GND nfet
M5 n2 g n1 GND nfet
M6 n3 h n2 GND nfet
M7 n3 i n2 GND nfet
M8 n3 j n2 GND nfet
M9 n3 b GND GND nfet
M10 n4 a n3 GND nfet
M11 n5 c VDD VDD pfet
M12 n4 d n5 VDD pfet
M13 n7 e VDD VDD pfet
M14 n8 f n7 VDD pfet
M15 n4 g n8 VDD pfet
M16 n10 h VDD VDD pfet
M17 n11 i n10 VDD pfet
M18 n4 j n11 VDD pfet
M19 n4 b n4 VDD pfet
M20 n4 a VDD VDD pfet
A equação é :(a*(b+(c+d+e)*(f+g+h)*(i+j+k)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n1 e GND GND nfet
M4 n2 f n1 GND nfet
M5 n2 g n1 GND nfet
M6 n2 h n1 GND nfet
M7 n3 i n2 GND nfet
M8 n3 j n2 GND nfet
M9 n3 k n2 GND nfet
M10 n3 b GND GND nfet
M11 n4 a n3 GND nfet
M12 n5 c VDD VDD pfet
M13 n6 d n5 VDD pfet
M14 n4 e n6 VDD pfet
M15 n8 f VDD VDD pfet
M16 n9 g n8 VDD pfet
M17 n4 h n9 VDD pfet
M18 n11 i VDD VDD pfet
M19 n12 j n11 VDD pfet
M20 n4 k n12 VDD pfet
M21 n4 b n4 VDD pfet
M22 n4 a VDD VDD pfet
A equação é :(a*(b*c+d*e))
M1 n1 b GND GND nfet
M2 n5 c n1 GND nfet
M3 n3 d GND GND nfet
M4 n5 e n3 GND nfet
M5 n5 a n5 GND nfet
M6 n6 b VDD VDD pfet
M7 n6 c VDD VDD pfet
M8 n5 d n6 VDD pfet
M9 n5 e n6 VDD pfet
M10 n5 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+f)))
M1 n1 b GND GND nfet
M2 n5 c n1 GND nfet
M3 n3 e GND GND nfet
M4 n3 f GND GND nfet
M5 n5 d n3 GND nfet
M6 n5 a n5 GND nfet
M7 n6 b VDD VDD pfet
M8 n6 c VDD VDD pfet
M9 n7 e n6 VDD pfet
M10 n5 f n7 VDD pfet
M11 n5 d n6 VDD pfet
M12 n5 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+f*g)))
M1 n1 b GND GND nfet
M2 n6 c n1 GND nfet
M3 n3 f GND GND nfet
M4 n4 g n3 GND nfet
M5 n4 e GND GND nfet
M6 n6 d n4 GND nfet
M7 n6 a n6 GND nfet
M8 n7 b VDD VDD pfet
M9 n7 c VDD VDD pfet
M10 n8 f n7 VDD pfet
M11 n8 g n7 VDD pfet
M12 n6 e n8 VDD pfet
M13 n6 d n7 VDD pfet
M14 n6 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+f*(g+h))))
M1 n1 b GND GND nfet
M2 n6 c n1 GND nfet
M3 n3 g GND GND nfet
M4 n3 h GND GND nfet
M5 n4 f n3 GND nfet
M6 n4 e GND GND nfet
M7 n6 d n4 GND nfet
M8 n6 a n6 GND nfet
M9 n7 b VDD VDD pfet
M10 n7 c VDD VDD pfet
M11 n8 g n7 VDD pfet
M12 n9 h n8 VDD pfet
M13 n9 f n7 VDD pfet
M14 n6 e n9 VDD pfet
M15 n6 d n7 VDD pfet
M16 n6 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+(f+g)*(h+i))))
M1 n1 b GND GND nfet
M2 n6 c n1 GND nfet
M3 n3 f GND GND nfet
M4 n3 g GND GND nfet
M5 n4 h n3 GND nfet
M6 n4 i n3 GND nfet
M7 n4 e GND GND nfet
M8 n6 d n4 GND nfet
M9 n6 a n6 GND nfet
M10 n7 b VDD VDD pfet
M11 n7 c VDD VDD pfet
M12 n8 f n7 VDD pfet
M13 n6 g n8 VDD pfet
M14 n10 h n7 VDD pfet
M15 n6 i n10 VDD pfet
M16 n6 e n6 VDD pfet
M17 n6 d n7 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b*c+d*(e*f+g*h)))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 e GND GND nfet
M4 n8 f n3 GND nfet
M5 n5 g GND GND nfet
M6 n8 h n5 GND nfet
M7 n8 d n8 GND nfet
M8 n8 a n8 GND nfet
M9 n9 b VDD VDD pfet
M10 n9 c VDD VDD pfet
M11 n10 e n9 VDD pfet
M12 n10 f n9 VDD pfet
M13 n8 g n10 VDD pfet
M14 n8 h n10 VDD pfet
M15 n8 d n9 VDD pfet
M16 n8 a VDD VDD pfet
A equação é :(a*(b*c+d*(e*f+g*(h+i))))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 e GND GND nfet
M4 n8 f n3 GND nfet
M5 n5 h GND GND nfet
M6 n5 i GND GND nfet
M7 n8 g n5 GND nfet
M8 n8 d n8 GND nfet
M9 n8 a n8 GND nfet
M10 n9 b VDD VDD pfet
M11 n9 c VDD VDD pfet
M12 n10 e n9 VDD pfet
M13 n10 f n9 VDD pfet
M14 n11 h n10 VDD pfet
M15 n8 i n11 VDD pfet
M16 n8 g n10 VDD pfet
M17 n8 d n9 VDD pfet
M18 n8 a VDD VDD pfet
A equação é :(a*(b*c+d*(e*f+(g+h)*(i+j))))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 g GND GND nfet
M4 n3 h GND GND nfet
M5 n8 i n3 GND nfet
M6 n8 j n3 GND nfet
M7 n5 e GND GND nfet
M8 n8 f n5 GND nfet
M9 n8 d n8 GND nfet
M10 n8 a n8 GND nfet
M11 n9 b VDD VDD pfet
M12 n9 c VDD VDD pfet
M13 n10 g n9 VDD pfet
M14 n8 h n10 VDD pfet
M15 n12 i n9 VDD pfet
M16 n8 j n12 VDD pfet
M17 n8 e n8 VDD pfet
M18 n8 f n8 VDD pfet
M19 n8 d n9 VDD pfet
M20 n8 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+f+g)))
M1 n1 b GND GND nfet
M2 n5 c n1 GND nfet
M3 n3 e GND GND nfet
M4 n3 f GND GND nfet
M5 n3 g GND GND nfet
M6 n5 d n3 GND nfet
M7 n5 a n5 GND nfet
M8 n6 b VDD VDD pfet
M9 n6 c VDD VDD pfet
M10 n7 e n6 VDD pfet
M11 n8 f n7 VDD pfet
M12 n5 g n8 VDD pfet
M13 n5 d n6 VDD pfet
M14 n5 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+f+g*h)))
M1 n1 b GND GND nfet
M2 n7 c n1 GND nfet
M3 n7 e GND GND nfet
M4 n7 f GND GND nfet
M5 n4 g GND GND nfet
M6 n7 h n4 GND nfet
M7 n7 d n7 GND nfet
M8 n7 a n7 GND nfet
M9 n8 b VDD VDD pfet
M10 n8 c VDD VDD pfet
M11 n9 e n8 VDD pfet
M12 n10 f n9 VDD pfet
M13 n7 g n10 VDD pfet
M14 n7 h n10 VDD pfet
M15 n7 d n8 VDD pfet
M16 n7 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+f*g+h*i)))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 f GND GND nfet
M4 n8 g n3 GND nfet
M5 n8 e GND GND nfet
M6 n5 h GND GND nfet
M7 n8 i n5 GND nfet
M8 n8 d n8 GND nfet
M9 n8 a n8 GND nfet
M10 n9 b VDD VDD pfet
M11 n9 c VDD VDD pfet
M12 n10 f n9 VDD pfet
M13 n10 g n9 VDD pfet
M14 n11 e n10 VDD pfet
M15 n8 h n11 VDD pfet
M16 n8 i n11 VDD pfet
M17 n8 d n9 VDD pfet
M18 n8 a VDD VDD pfet
A equação é :(a*(b*c+d*(e*f+g*h+i*j)))
M1 n1 b GND GND nfet
M2 n10 c n1 GND nfet
M3 n3 e GND GND nfet
M4 n10 f n3 GND nfet
M5 n5 g GND GND nfet
M6 n10 h n5 GND nfet
M7 n7 i GND GND nfet
M8 n10 j n7 GND nfet
M9 n10 d n10 GND nfet
M10 n10 a n10 GND nfet
M11 n11 b VDD VDD pfet
M12 n11 c VDD VDD pfet
M13 n12 e n11 VDD pfet
M14 n12 f n11 VDD pfet
M15 n13 g n12 VDD pfet
M16 n13 h n12 VDD pfet
M17 n10 i n13 VDD pfet
M18 n10 j n13 VDD pfet
M19 n10 d n11 VDD pfet
M20 n10 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+g)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n5 f n1 GND nfet
M4 n5 g n1 GND nfet
M5 n3 b GND GND nfet
M6 n5 c n3 GND nfet
M7 n5 a n5 GND nfet
M8 n6 d VDD VDD pfet
M9 n5 e n6 VDD pfet
M10 n8 f VDD VDD pfet
M11 n5 g n8 VDD pfet
M12 n5 b n5 VDD pfet
M13 n5 c n5 VDD pfet
M14 n5 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+g*h)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n2 g n1 GND nfet
M4 n6 h n2 GND nfet
M5 n6 f n1 GND nfet
M6 n4 b GND GND nfet
M7 n6 c n4 GND nfet
M8 n6 a n6 GND nfet
M9 n7 d VDD VDD pfet
M10 n6 e n7 VDD pfet
M11 n9 g VDD VDD pfet
M12 n9 h VDD VDD pfet
M13 n6 f n9 VDD pfet
M14 n6 b n6 VDD pfet
M15 n6 c n6 VDD pfet
M16 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+g*(h+i))))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n2 h n1 GND nfet
M4 n2 i n1 GND nfet
M5 n6 g n2 GND nfet
M6 n6 f n1 GND nfet
M7 n4 b GND GND nfet
M8 n6 c n4 GND nfet
M9 n6 a n6 GND nfet
M10 n7 d VDD VDD pfet
M11 n6 e n7 VDD pfet
M12 n9 h VDD VDD pfet
M13 n10 i n9 VDD pfet
M14 n10 g VDD VDD pfet
M15 n6 f n10 VDD pfet
M16 n6 b n6 VDD pfet
M17 n6 c n6 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+(g+h)*(i+j))))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n6 i n2 GND nfet
M6 n6 j n2 GND nfet
M7 n6 f n1 GND nfet
M8 n4 b GND GND nfet
M9 n6 c n4 GND nfet
M10 n6 a n6 GND nfet
M11 n7 d VDD VDD pfet
M12 n6 e n7 VDD pfet
M13 n9 g VDD VDD pfet
M14 n6 h n9 VDD pfet
M15 n11 i VDD VDD pfet
M16 n6 j n11 VDD pfet
M17 n6 f n6 VDD pfet
M18 n6 b n6 VDD pfet
M19 n6 c n6 VDD pfet
M20 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f*g+h*i)))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 f GND GND nfet
M4 n8 g n3 GND nfet
M5 n5 h GND GND nfet
M6 n8 i n5 GND nfet
M7 n8 d n8 GND nfet
M8 n8 e n8 GND nfet
M9 n8 a n8 GND nfet
M10 n9 b VDD VDD pfet
M11 n9 c VDD VDD pfet
M12 n10 f n9 VDD pfet
M13 n10 g n9 VDD pfet
M14 n8 h n10 VDD pfet
M15 n8 i n10 VDD pfet
M16 n12 d n9 VDD pfet
M17 n8 e n12 VDD pfet
M18 n8 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f*g+h*(i+j))))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 f GND GND nfet
M4 n8 g n3 GND nfet
M5 n5 i GND GND nfet
M6 n5 j GND GND nfet
M7 n8 h n5 GND nfet
M8 n8 d n8 GND nfet
M9 n8 e n8 GND nfet
M10 n8 a n8 GND nfet
M11 n9 b VDD VDD pfet
M12 n9 c VDD VDD pfet
M13 n10 f n9 VDD pfet
M14 n10 g n9 VDD pfet
M15 n11 i n10 VDD pfet
M16 n8 j n11 VDD pfet
M17 n8 h n10 VDD pfet
M18 n13 d n9 VDD pfet
M19 n8 e n13 VDD pfet
M20 n8 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f*g+(h+i)*(j+k))))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n2 h n1 GND nfet
M4 n2 i n1 GND nfet
M5 n8 j n2 GND nfet
M6 n8 k n2 GND nfet
M7 n4 f n1 GND nfet
M8 n8 g n4 GND nfet
M9 n6 b GND GND nfet
M10 n8 c n6 GND nfet
M11 n8 a n8 GND nfet
M12 n9 d VDD VDD pfet
M13 n8 e n9 VDD pfet
M14 n11 h VDD VDD pfet
M15 n8 i n11 VDD pfet
M16 n13 j VDD VDD pfet
M17 n8 k n13 VDD pfet
M18 n8 f n8 VDD pfet
M19 n8 g n8 VDD pfet
M20 n8 b n8 VDD pfet
M21 n8 c n8 VDD pfet
M22 n8 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+g+h)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n5 f n1 GND nfet
M4 n5 g n1 GND nfet
M5 n5 h n1 GND nfet
M6 n3 b GND GND nfet
M7 n5 c n3 GND nfet
M8 n5 a n5 GND nfet
M9 n6 d VDD VDD pfet
M10 n5 e n6 VDD pfet
M11 n8 f VDD VDD pfet
M12 n9 g n8 VDD pfet
M13 n5 h n9 VDD pfet
M14 n5 b n5 VDD pfet
M15 n5 c n5 VDD pfet
M16 n5 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+g+h*i)))
M1 n1 b GND GND nfet
M2 n7 c n1 GND nfet
M3 n7 f GND GND nfet
M4 n7 g GND GND nfet
M5 n4 h GND GND nfet
M6 n7 i n4 GND nfet
M7 n7 d n7 GND nfet
M8 n7 e n7 GND nfet
M9 n7 a n7 GND nfet
M10 n8 b VDD VDD pfet
M11 n8 c VDD VDD pfet
M12 n9 f n8 VDD pfet
M13 n10 g n9 VDD pfet
M14 n7 h n10 VDD pfet
M15 n7 i n10 VDD pfet
M16 n12 d n8 VDD pfet
M17 n7 e n12 VDD pfet
M18 n7 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+g*h+i*j)))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 g GND GND nfet
M4 n8 h n3 GND nfet
M5 n8 f GND GND nfet
M6 n5 i GND GND nfet
M7 n8 j n5 GND nfet
M8 n8 d n8 GND nfet
M9 n8 e n8 GND nfet
M10 n8 a n8 GND nfet
M11 n9 b VDD VDD pfet
M12 n9 c VDD VDD pfet
M13 n10 g n9 VDD pfet
M14 n10 h n9 VDD pfet
M15 n11 f n10 VDD pfet
M16 n8 i n11 VDD pfet
M17 n8 j n11 VDD pfet
M18 n13 d n9 VDD pfet
M19 n8 e n13 VDD pfet
M20 n8 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f*g+h*i+j*k)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n2 f n1 GND nfet
M4 n10 g n2 GND nfet
M5 n4 h n1 GND nfet
M6 n10 i n4 GND nfet
M7 n6 j n1 GND nfet
M8 n10 k n6 GND nfet
M9 n8 b GND GND nfet
M10 n10 c n8 GND nfet
M11 n10 a n10 GND nfet
M12 n11 d VDD VDD pfet
M13 n10 e n11 VDD pfet
M14 n13 f VDD VDD pfet
M15 n13 g VDD VDD pfet
M16 n14 h n13 VDD pfet
M17 n14 i n13 VDD pfet
M18 n10 j n14 VDD pfet
M19 n10 k n14 VDD pfet
M20 n10 b n10 VDD pfet
M21 n10 c n10 VDD pfet
M22 n10 a VDD VDD pfet
A equação é :(a*(b*c+(d+e*f)*(g+h+i)))
M1 n1 e GND GND nfet
M2 n2 f n1 GND nfet
M3 n2 d GND GND nfet
M4 n6 g n2 GND nfet
M5 n6 h n2 GND nfet
M6 n6 i n2 GND nfet
M7 n4 b GND GND nfet
M8 n6 c n4 GND nfet
M9 n6 a n6 GND nfet
M10 n7 e VDD VDD pfet
M11 n7 f VDD VDD pfet
M12 n6 d n7 VDD pfet
M13 n9 g VDD VDD pfet
M14 n10 h n9 VDD pfet
M15 n6 i n10 VDD pfet
M16 n6 b n6 VDD pfet
M17 n6 c n6 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d+e*(f+g))*(h+i+j)))
M1 n1 f GND GND nfet
M2 n1 g GND GND nfet
M3 n2 e n1 GND nfet
M4 n2 d GND GND nfet
M5 n6 h n2 GND nfet
M6 n6 i n2 GND nfet
M7 n6 j n2 GND nfet
M8 n4 b GND GND nfet
M9 n6 c n4 GND nfet
M10 n6 a n6 GND nfet
M11 n7 f VDD VDD pfet
M12 n8 g n7 VDD pfet
M13 n8 e VDD VDD pfet
M14 n6 d n8 VDD pfet
M15 n10 h VDD VDD pfet
M16 n11 i n10 VDD pfet
M17 n6 j n11 VDD pfet
M18 n6 b n6 VDD pfet
M19 n6 c n6 VDD pfet
M20 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d+(e+f)*(g+h))*(i+j+k)))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 g n1 GND nfet
M4 n2 h n1 GND nfet
M5 n2 d GND GND nfet
M6 n6 i n2 GND nfet
M7 n6 j n2 GND nfet
M8 n6 k n2 GND nfet
M9 n4 b GND GND nfet
M10 n6 c n4 GND nfet
M11 n6 a n6 GND nfet
M12 n7 e VDD VDD pfet
M13 n6 f n7 VDD pfet
M14 n9 g VDD VDD pfet
M15 n6 h n9 VDD pfet
M16 n6 d n6 VDD pfet
M17 n12 i VDD VDD pfet
M18 n13 j n12 VDD pfet
M19 n6 k n13 VDD pfet
M20 n6 b n6 VDD pfet
M21 n6 c n6 VDD pfet
M22 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d*e+f*g)*(h+i+j)))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 d GND GND nfet
M4 n8 e n3 GND nfet
M5 n5 f GND GND nfet
M6 n8 g n5 GND nfet
M7 n8 h n8 GND nfet
M8 n8 i n8 GND nfet
M9 n8 j n8 GND nfet
M10 n8 a n8 GND nfet
M11 n9 b VDD VDD pfet
M12 n9 c VDD VDD pfet
M13 n10 d n9 VDD pfet
M14 n10 e n9 VDD pfet
M15 n8 f n10 VDD pfet
M16 n8 g n10 VDD pfet
M17 n12 h n9 VDD pfet
M18 n13 i n12 VDD pfet
M19 n8 j n13 VDD pfet
M20 n8 a VDD VDD pfet
A equação é :(a*(b*c+(d*e+f*(g+h))*(i+j+k)))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 d GND GND nfet
M4 n8 e n3 GND nfet
M5 n5 g GND GND nfet
M6 n5 h GND GND nfet
M7 n8 f n5 GND nfet
M8 n8 i n8 GND nfet
M9 n8 j n8 GND nfet
M10 n8 k n8 GND nfet
M11 n8 a n8 GND nfet
M12 n9 b VDD VDD pfet
M13 n9 c VDD VDD pfet
M14 n10 d n9 VDD pfet
M15 n10 e n9 VDD pfet
M16 n11 g n10 VDD pfet
M17 n8 h n11 VDD pfet
M18 n8 f n10 VDD pfet
M19 n13 i n9 VDD pfet
M20 n14 j n13 VDD pfet
M21 n8 k n14 VDD pfet
M22 n8 a VDD VDD pfet
A equação é :(a*(b*c+(d*e+(f+g)*(h+i))*(j+k+l)))
M1 n1 f GND GND nfet
M2 n1 g GND GND nfet
M3 n8 h n1 GND nfet
M4 n8 i n1 GND nfet
M5 n3 d GND GND nfet
M6 n8 e n3 GND nfet
M7 n8 j n8 GND nfet
M8 n8 k n8 GND nfet
M9 n8 l n8 GND nfet
M10 n6 b GND GND nfet
M11 n8 c n6 GND nfet
M12 n8 a n8 GND nfet
M13 n9 f VDD VDD pfet
M14 n8 g n9 VDD pfet
M15 n11 h VDD VDD pfet
M16 n8 i n11 VDD pfet
M17 n8 d n8 VDD pfet
M18 n8 e n8 VDD pfet
M19 n14 j VDD VDD pfet
M20 n15 k n14 VDD pfet
M21 n8 l n15 VDD pfet
M22 n8 b n8 VDD pfet
M23 n8 c n8 VDD pfet
M24 n8 a VDD VDD pfet
A equação é :(a*(b*c+(d+e+f)*(g+h+i)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n1 f GND GND nfet
M4 n5 g n1 GND nfet
M5 n5 h n1 GND nfet
M6 n5 i n1 GND nfet
M7 n3 b GND GND nfet
M8 n5 c n3 GND nfet
M9 n5 a n5 GND nfet
M10 n6 d VDD VDD pfet
M11 n7 e n6 VDD pfet
M12 n5 f n7 VDD pfet
M13 n9 g VDD VDD pfet
M14 n10 h n9 VDD pfet
M15 n5 i n10 VDD pfet
M16 n5 b n5 VDD pfet
M17 n5 c n5 VDD pfet
M18 n5 a VDD VDD pfet
A equação é :(a*(b*c+(d+e+f)*(g+h+i*j)))
M1 n1 b GND GND nfet
M2 n7 c n1 GND nfet
M3 n7 g GND GND nfet
M4 n7 h GND GND nfet
M5 n4 i GND GND nfet
M6 n7 j n4 GND nfet
M7 n7 d n7 GND nfet
M8 n7 e n7 GND nfet
M9 n7 f n7 GND nfet
M10 n7 a n7 GND nfet
M11 n8 b VDD VDD pfet
M12 n8 c VDD VDD pfet
M13 n9 g n8 VDD pfet
M14 n10 h n9 VDD pfet
M15 n7 i n10 VDD pfet
M16 n7 j n10 VDD pfet
M17 n12 d n8 VDD pfet
M18 n13 e n12 VDD pfet
M19 n7 f n13 VDD pfet
M20 n7 a VDD VDD pfet
A equação é :(a*(b*c+(d+e+f)*(g+h*i+j*k)))
M1 n1 b GND GND nfet
M2 n8 c n1 GND nfet
M3 n3 h GND GND nfet
M4 n8 i n3 GND nfet
M5 n8 g GND GND nfet
M6 n5 j GND GND nfet
M7 n8 k n5 GND nfet
M8 n8 d n8 GND nfet
M9 n8 e n8 GND nfet
M10 n8 f n8 GND nfet
M11 n8 a n8 GND nfet
M12 n9 b VDD VDD pfet
M13 n9 c VDD VDD pfet
M14 n10 h n9 VDD pfet
M15 n10 i n9 VDD pfet
M16 n11 g n10 VDD pfet
M17 n8 j n11 VDD pfet
M18 n8 k n11 VDD pfet
M19 n13 d n9 VDD pfet
M20 n14 e n13 VDD pfet
M21 n8 f n14 VDD pfet
M22 n8 a VDD VDD pfet
A equação é :(a*(b*c+(d+e+f)*(g*h+i*j+k*l)))
M1 n1 d GND GND nfet
M2 n1 e GND GND nfet
M3 n1 f GND GND nfet
M4 n2 g n1 GND nfet
M5 n10 h n2 GND nfet
M6 n4 i n1 GND nfet
M7 n10 j n4 GND nfet
M8 n6 k n1 GND nfet
M9 n10 l n6 GND nfet
M10 n8 b GND GND nfet
M11 n10 c n8 GND nfet
M12 n10 a n10 GND nfet
M13 n11 d VDD VDD pfet
M14 n12 e n11 VDD pfet
M15 n10 f n12 VDD pfet
M16 n14 g VDD VDD pfet
M17 n14 h VDD VDD pfet
M18 n15 i n14 VDD pfet
M19 n15 j n14 VDD pfet
M20 n10 k n15 VDD pfet
M21 n10 l n15 VDD pfet
M22 n10 b n10 VDD pfet
M23 n10 c n10 VDD pfet
M24 n10 a VDD VDD pfet
A equação é :(a*(b*c+d*e*f))
M1 n1 b GND GND nfet
M2 n6 c n1 GND nfet
M3 n3 d GND GND nfet
M4 n4 e n3 GND nfet
M5 n6 f n4 GND nfet
M6 n6 a n6 GND nfet
M7 n7 b VDD VDD pfet
M8 n7 c VDD VDD pfet
M9 n6 d n7 VDD pfet
M10 n6 e n7 VDD pfet
M11 n6 f n7 VDD pfet
M12 n6 a VDD VDD pfet
A equação é :(a*(b*c+d*e*(f+g)))
M1 n1 d GND GND nfet
M2 n2 e n1 GND nfet
M3 n6 f n2 GND nfet
M4 n6 g n2 GND nfet
M5 n4 b GND GND nfet
M6 n6 c n4 GND nfet
M7 n6 a n6 GND nfet
M8 n6 d VDD VDD pfet
M9 n6 e VDD VDD pfet
M10 n8 f VDD VDD pfet
M11 n6 g n8 VDD pfet
M12 n6 b n6 VDD pfet
M13 n6 c n6 VDD pfet
M14 n6 a VDD VDD pfet
A equação é :(a*(b*c+d*e*(f+g+h)))
M1 n1 d GND GND nfet
M2 n2 e n1 GND nfet
M3 n6 f n2 GND nfet
M4 n6 g n2 GND nfet
M5 n6 h n2 GND nfet
M6 n4 b GND GND nfet
M7 n6 c n4 GND nfet
M8 n6 a n6 GND nfet
M9 n6 d VDD VDD pfet
M10 n6 e VDD VDD pfet
M11 n8 f VDD VDD pfet
M12 n9 g n8 VDD pfet
M13 n6 h n9 VDD pfet
M14 n6 b n6 VDD pfet
M15 n6 c n6 VDD pfet
M16 n6 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+f)*(g+h)))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 d n1 GND nfet
M4 n6 g n2 GND nfet
M5 n6 h n2 GND nfet
M6 n4 b GND GND nfet
M7 n6 c n4 GND nfet
M8 n6 a n6 GND nfet
M9 n7 e VDD VDD pfet
M10 n6 f n7 VDD pfet
M11 n6 d VDD VDD pfet
M12 n9 g VDD VDD pfet
M13 n6 h n9 VDD pfet
M14 n6 b n6 VDD pfet
M15 n6 c n6 VDD pfet
M16 n6 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+f)*(g+h+i)))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 d n1 GND nfet
M4 n6 g n2 GND nfet
M5 n6 h n2 GND nfet
M6 n6 i n2 GND nfet
M7 n4 b GND GND nfet
M8 n6 c n4 GND nfet
M9 n6 a n6 GND nfet
M10 n7 e VDD VDD pfet
M11 n6 f n7 VDD pfet
M12 n6 d VDD VDD pfet
M13 n9 g VDD VDD pfet
M14 n10 h n9 VDD pfet
M15 n6 i n10 VDD pfet
M16 n6 b n6 VDD pfet
M17 n6 c n6 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b*c+d*(e+f+g)*(h+i+j)))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n1 g GND GND nfet
M4 n2 d n1 GND nfet
M5 n6 h n2 GND nfet
M6 n6 i n2 GND nfet
M7 n6 j n2 GND nfet
M8 n4 b GND GND nfet
M9 n6 c n4 GND nfet
M10 n6 a n6 GND nfet
M11 n7 e VDD VDD pfet
M12 n8 f n7 VDD pfet
M13 n6 g n8 VDD pfet
M14 n6 d VDD VDD pfet
M15 n10 h VDD VDD pfet
M16 n11 i n10 VDD pfet
M17 n6 j n11 VDD pfet
M18 n6 b n6 VDD pfet
M19 n6 c n6 VDD pfet
M20 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+g)*(h+i)))
M1 n1 b GND GND nfet
M2 n6 c n1 GND nfet
M3 n3 d GND GND nfet
M4 n3 e GND GND nfet
M5 n4 f n3 GND nfet
M6 n4 g n3 GND nfet
M7 n6 h n4 GND nfet
M8 n6 i n4 GND nfet
M9 n6 a n6 GND nfet
M10 n7 b VDD VDD pfet
M11 n7 c VDD VDD pfet
M12 n8 d n7 VDD pfet
M13 n6 e n8 VDD pfet
M14 n10 f n7 VDD pfet
M15 n6 g n10 VDD pfet
M16 n12 h n7 VDD pfet
M17 n6 i n12 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+g)*(h+i+j)))
M1 n1 b GND GND nfet
M2 n6 c n1 GND nfet
M3 n3 d GND GND nfet
M4 n3 e GND GND nfet
M5 n4 f n3 GND nfet
M6 n4 g n3 GND nfet
M7 n6 h n4 GND nfet
M8 n6 i n4 GND nfet
M9 n6 j n4 GND nfet
M10 n6 a n6 GND nfet
M11 n7 b VDD VDD pfet
M12 n7 c VDD VDD pfet
M13 n8 d n7 VDD pfet
M14 n6 e n8 VDD pfet
M15 n10 f n7 VDD pfet
M16 n6 g n10 VDD pfet
M17 n12 h n7 VDD pfet
M18 n13 i n12 VDD pfet
M19 n6 j n13 VDD pfet
M20 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d+e)*(f+g+h)*(i+j+k)))
M1 n1 b GND GND nfet
M2 n6 c n1 GND nfet
M3 n3 d GND GND nfet
M4 n3 e GND GND nfet
M5 n4 f n3 GND nfet
M6 n4 g n3 GND nfet
M7 n4 h n3 GND nfet
M8 n6 i n4 GND nfet
M9 n6 j n4 GND nfet
M10 n6 k n4 GND nfet
M11 n6 a n6 GND nfet
M12 n7 b VDD VDD pfet
M13 n7 c VDD VDD pfet
M14 n8 d n7 VDD pfet
M15 n6 e n8 VDD pfet
M16 n10 f n7 VDD pfet
M17 n11 g n10 VDD pfet
M18 n6 h n11 VDD pfet
M19 n13 i n7 VDD pfet
M20 n14 j n13 VDD pfet
M21 n6 k n14 VDD pfet
M22 n6 a VDD VDD pfet
A equação é :(a*(b*c+(d+e+f)*(g+h+i)*(j+k+l)))
M1 n1 b GND GND nfet
M2 n6 c n1 GND nfet
M3 n3 d GND GND nfet
M4 n3 e GND GND nfet
M5 n3 f GND GND nfet
M6 n4 g n3 GND nfet
M7 n4 h n3 GND nfet
M8 n4 i n3 GND nfet
M9 n6 j n4 GND nfet
M10 n6 k n4 GND nfet
M11 n6 l n4 GND nfet
M12 n6 a n6 GND nfet
M13 n7 b VDD VDD pfet
M14 n7 c VDD VDD pfet
M15 n8 d n7 VDD pfet
M16 n9 e n8 VDD pfet
M17 n6 f n9 VDD pfet
M18 n11 g n7 VDD pfet
M19 n12 h n11 VDD pfet
M20 n6 i n12 VDD pfet
M21 n14 j n7 VDD pfet
M22 n15 k n14 VDD pfet
M23 n6 l n15 VDD pfet
M24 n6 a VDD VDD pfet
A equação é :(a*(b*(c+d)+e*(f+g)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n5 b n1 GND nfet
M4 n3 f GND GND nfet
M5 n3 g GND GND nfet
M6 n5 e n3 GND nfet
M7 n5 a n5 GND nfet
M8 n6 c VDD VDD pfet
M9 n7 d n6 VDD pfet
M10 n7 b VDD VDD pfet
M11 n8 f n7 VDD pfet
M12 n5 g n8 VDD pfet
M13 n5 e n7 VDD pfet
M14 n5 a VDD VDD pfet
A equação é :(a*(b*(c+d)+e*(f+g*h)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n6 b n1 GND nfet
M4 n3 g GND GND nfet
M5 n4 h n3 GND nfet
M6 n4 f GND GND nfet
M7 n6 e n4 GND nfet
M8 n6 a n6 GND nfet
M9 n7 c VDD VDD pfet
M10 n8 d n7 VDD pfet
M11 n8 b VDD VDD pfet
M12 n9 g n8 VDD pfet
M13 n9 h n8 VDD pfet
M14 n6 f n9 VDD pfet
M15 n6 e n8 VDD pfet
M16 n6 a VDD VDD pfet
A equação é :(a*(b*(c+d)+e*(f*g+h*i)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n8 b n1 GND nfet
M4 n3 f GND GND nfet
M5 n8 g n3 GND nfet
M6 n5 h GND GND nfet
M7 n8 i n5 GND nfet
M8 n8 e n8 GND nfet
M9 n8 a n8 GND nfet
M10 n9 c VDD VDD pfet
M11 n10 d n9 VDD pfet
M12 n10 b VDD VDD pfet
M13 n11 f n10 VDD pfet
M14 n11 g n10 VDD pfet
M15 n8 h n11 VDD pfet
M16 n8 i n11 VDD pfet
M17 n8 e n10 VDD pfet
M18 n8 a VDD VDD pfet
A equação é :(a*(b*(c+d)+(e+f)*(g+h)))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n5 g n1 GND nfet
M4 n5 h n1 GND nfet
M5 n3 c GND GND nfet
M6 n3 d GND GND nfet
M7 n5 b n3 GND nfet
M8 n5 a n5 GND nfet
M9 n6 e VDD VDD pfet
M10 n5 f n6 VDD pfet
M11 n8 g VDD VDD pfet
M12 n5 h n8 VDD pfet
M13 n10 c n5 VDD pfet
M14 n5 d n10 VDD pfet
M15 n5 b n5 VDD pfet
M16 n5 a VDD VDD pfet
A equação é :(a*(b*(c+d)+(e+f)*(g+h*i)))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 h n1 GND nfet
M4 n6 i n2 GND nfet
M5 n6 g n1 GND nfet
M6 n4 c GND GND nfet
M7 n4 d GND GND nfet
M8 n6 b n4 GND nfet
M9 n6 a n6 GND nfet
M10 n7 e VDD VDD pfet
M11 n6 f n7 VDD pfet
M12 n9 h VDD VDD pfet
M13 n9 i VDD VDD pfet
M14 n6 g n9 VDD pfet
M15 n11 c n6 VDD pfet
M16 n6 d n11 VDD pfet
M17 n6 b n6 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b*(c+d)+(e+f)*(g*h+i*j)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n8 b n1 GND nfet
M4 n3 g GND GND nfet
M5 n8 h n3 GND nfet
M6 n5 i GND GND nfet
M7 n8 j n5 GND nfet
M8 n8 e n8 GND nfet
M9 n8 f n8 GND nfet
M10 n8 a n8 GND nfet
M11 n9 c VDD VDD pfet
M12 n10 d n9 VDD pfet
M13 n10 b VDD VDD pfet
M14 n11 g n10 VDD pfet
M15 n11 h n10 VDD pfet
M16 n8 i n11 VDD pfet
M17 n8 j n11 VDD pfet
M18 n13 e n10 VDD pfet
M19 n8 f n13 VDD pfet
M20 n8 a VDD VDD pfet
A equação é :(a*(b*(c+d)+e*f*g))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n6 b n1 GND nfet
M4 n3 e GND GND nfet
M5 n4 f n3 GND nfet
M6 n6 g n4 GND nfet
M7 n6 a n6 GND nfet
M8 n7 c VDD VDD pfet
M9 n8 d n7 VDD pfet
M10 n8 b VDD VDD pfet
M11 n6 e n8 VDD pfet
M12 n6 f n8 VDD pfet
M13 n6 g n8 VDD pfet
M14 n6 a VDD VDD pfet
A equação é :(a*(b*(c+d)+e*f*(g+h)))
M1 n1 e GND GND nfet
M2 n2 f n1 GND nfet
M3 n6 g n2 GND nfet
M4 n6 h n2 GND nfet
M5 n4 c GND GND nfet
M6 n4 d GND GND nfet
M7 n6 b n4 GND nfet
M8 n6 a n6 GND nfet
M9 n6 e VDD VDD pfet
M10 n6 f VDD VDD pfet
M11 n8 g VDD VDD pfet
M12 n6 h n8 VDD pfet
M13 n10 c n6 VDD pfet
M14 n6 d n10 VDD pfet
M15 n6 b n6 VDD pfet
M16 n6 a VDD VDD pfet
A equação é :(a*(b*(c+d)+e*(f+g)*(h+i)))
M1 n1 f GND GND nfet
M2 n1 g GND GND nfet
M3 n2 e n1 GND nfet
M4 n6 h n2 GND nfet
M5 n6 i n2 GND nfet
M6 n4 c GND GND nfet
M7 n4 d GND GND nfet
M8 n6 b n4 GND nfet
M9 n6 a n6 GND nfet
M10 n7 f VDD VDD pfet
M11 n6 g n7 VDD pfet
M12 n6 e VDD VDD pfet
M13 n9 h VDD VDD pfet
M14 n6 i n9 VDD pfet
M15 n11 c n6 VDD pfet
M16 n6 d n11 VDD pfet
M17 n6 b n6 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b*(c+d)+(e+f)*(g+h)*(i+j)))
M1 n1 c GND GND nfet
M2 n1 d GND GND nfet
M3 n6 b n1 GND nfet
M4 n3 e GND GND nfet
M5 n3 f GND GND nfet
M6 n4 g n3 GND nfet
M7 n4 h n3 GND nfet
M8 n6 i n4 GND nfet
M9 n6 j n4 GND nfet
M10 n6 a n6 GND nfet
M11 n7 c VDD VDD pfet
M12 n8 d n7 VDD pfet
M13 n8 b VDD VDD pfet
M14 n9 e n8 VDD pfet
M15 n6 f n9 VDD pfet
M16 n11 g n8 VDD pfet
M17 n6 h n11 VDD pfet
M18 n13 i n8 VDD pfet
M19 n6 j n13 VDD pfet
M20 n6 a VDD VDD pfet
A equação é :(a*(b*(c+d*e)+f*(g+h*i)))
M1 n1 d GND GND nfet
M2 n2 e n1 GND nfet
M3 n2 c GND GND nfet
M4 n7 b n2 GND nfet
M5 n4 h GND GND nfet
M6 n5 i n4 GND nfet
M7 n5 g GND GND nfet
M8 n7 f n5 GND nfet
M9 n7 a n7 GND nfet
M10 n8 d VDD VDD pfet
M11 n8 e VDD VDD pfet
M12 n9 c n8 VDD pfet
M13 n9 b VDD VDD pfet
M14 n10 h n9 VDD pfet
M15 n10 i n9 VDD pfet
M16 n7 g n10 VDD pfet
M17 n7 f n9 VDD pfet
M18 n7 a VDD VDD pfet
A equação é :(a*(b*(c+d*e)+f*(g*h+i*j)))
M1 n1 d GND GND nfet
M2 n2 e n1 GND nfet
M3 n2 c GND GND nfet
M4 n9 b n2 GND nfet
M5 n4 g GND GND nfet
M6 n9 h n4 GND nfet
M7 n6 i GND GND nfet
M8 n9 j n6 GND nfet
M9 n9 f n9 GND nfet
M10 n9 a n9 GND nfet
M11 n10 d VDD VDD pfet
M12 n10 e VDD VDD pfet
M13 n11 c n10 VDD pfet
M14 n11 b VDD VDD pfet
M15 n12 g n11 VDD pfet
M16 n12 h n11 VDD pfet
M17 n9 i n12 VDD pfet
M18 n9 j n12 VDD pfet
M19 n9 f n11 VDD pfet
M20 n9 a VDD VDD pfet
A equação é :(a*(b*(c+d*e)+(f+g)*(h+i)))
M1 n1 f GND GND nfet
M2 n1 g GND GND nfet
M3 n6 h n1 GND nfet
M4 n6 i n1 GND nfet
M5 n3 d GND GND nfet
M6 n4 e n3 GND nfet
M7 n4 c GND GND nfet
M8 n6 b n4 GND nfet
M9 n6 a n6 GND nfet
M10 n7 f VDD VDD pfet
M11 n6 g n7 VDD pfet
M12 n9 h VDD VDD pfet
M13 n6 i n9 VDD pfet
M14 n11 d n6 VDD pfet
M15 n11 e n6 VDD pfet
M16 n6 c n11 VDD pfet
M17 n6 b n6 VDD pfet
M18 n6 a VDD VDD pfet
A equação é :(a*(b*(c+d*e)+(f+g)*(h+i*j)))
M1 n1 f GND GND nfet
M2 n1 g GND GND nfet
M3 n2 i n1 GND nfet
M4 n7 j n2 GND nfet
M5 n7 h n1 GND nfet
M6 n4 d GND GND nfet
M7 n5 e n4 GND nfet
M8 n5 c GND GND nfet
M9 n7 b n5 GND nfet
M10 n7 a n7 GND nfet
M11 n8 f VDD VDD pfet
M12 n7 g n8 VDD pfet
M13 n10 i VDD VDD pfet
M14 n10 j VDD VDD pfet
M15 n7 h n10 VDD pfet
M16 n12 d n7 VDD pfet
M17 n12 e n7 VDD pfet
M18 n7 c n12 VDD pfet
M19 n7 b n7 VDD pfet
M20 n7 a VDD VDD pfet
A equação é :(a*(b*(c+d*e)+(f+g)*(h*i+j*k)))
M1 n1 d GND GND nfet
M2 n2 e n1 GND nfet
M3 n2 c GND GND nfet
M4 n9 b n2 GND nfet
M5 n4 h GND GND nfet
M6 n9 i n4 GND nfet
M7 n6 j GND GND nfet
M8 n9 k n6 GND nfet
M9 n9 f n9 GND nfet
M10 n9 g n9 GND nfet
M11 n9 a n9 GND nfet
M12 n10 d VDD VDD pfet
M13 n10 e VDD VDD pfet
M14 n11 c n10 VDD pfet
M15 n11 b VDD VDD pfet
M16 n12 h n11 VDD pfet
M17 n12 i n11 VDD pfet
M18 n9 j n12 VDD pfet
M19 n9 k n12 VDD pfet
M20 n14 f n11 VDD pfet
M21 n9 g n14 VDD pfet
M22 n9 a VDD VDD pfet
A equação é :(a*(b*(c+d*e)+f*g*h))
M1 n1 d GND GND nfet
M2 n2 e n1 GND nfet
M3 n2 c GND GND nfet
M4 n7 b n2 GND nfet
M5 n4 f GND GND nfet
M6 n5 g n4 GND nfet
M7 n7 h n5 GND nfet
M8 n7 a n7 GND nfet
M9 n8 d VDD VDD pfet
M10 n8 e VDD VDD pfet
M11 n9 c n8 VDD pfet
M12 n9 b VDD VDD pfet
M13 n7 f n9 VDD pfet
M14 n7 g n9 VDD pfet
M15 n7 h n9 VDD pfet
M16 n7 a VDD VDD pfet
A equação é :(a*(b*(c+d*e)+f*g*(h+i)))
M1 n1 f GND GND nfet
M2 n2 g n1 GND nfet
M3 n7 h n2 GND nfet
M4 n7 i n2 GND nfet
M5 n4 d GND GND nfet
M6 n5 e n4 GND nfet
M7 n5 c GND GND nfet
M8 n7 b n5 GND nfet
M9 n7 a n7 GND nfet
M10 n7 f VDD VDD pfet
M11 n7 g VDD VDD pfet
M12 n9 h VDD VDD pfet
M13 n7 i n9 VDD pfet
M14 n11 d n7 VDD pfet
M15 n11 e n7 VDD pfet
M16 n7 c n11 VDD pfet
M17 n7 b n7 VDD pfet
M18 n7 a VDD VDD pfet
A equação é :(a*(b*(c+d*e)+f*(g+h)*(i+j)))
M1 n1 g GND GND nfet
M2 n1 h GND GND nfet
M3 n2 f n1 GND nfet
M4 n7 i n2 GND nfet
M5 n7 j n2 GND nfet
M6 n4 d GND GND nfet
M7 n5 e n4 GND nfet
M8 n5 c GND GND nfet
M9 n7 b n5 GND nfet
M10 n7 a n7 GND nfet
M11 n8 g VDD VDD pfet
M12 n7 h n8 VDD pfet
M13 n7 f VDD VDD pfet
M14 n10 i VDD VDD pfet
M15 n7 j n10 VDD pfet
M16 n12 d n7 VDD pfet
M17 n12 e n7 VDD pfet
M18 n7 c n12 VDD pfet
M19 n7 b n7 VDD pfet
M20 n7 a VDD VDD pfet
A equação é :(a*(b*(c+d*e)+(f+g)*(h+i)*(j+k)))
M1 n1 d GND GND nfet
M2 n2 e n1 GND nfet
M3 n2 c GND GND nfet
M4 n7 b n2 GND nfet
M5 n4 f GND GND nfet
M6 n4 g GND GND nfet
M7 n5 h n4 GND nfet
M8 n5 i n4 GND nfet
M9 n7 j n5 GND nfet
M10 n7 k n5 GND nfet
M11 n7 a n7 GND nfet
M12 n8 d VDD VDD pfet
M13 n8 e VDD VDD pfet
M14 n9 c n8 VDD pfet
M15 n9 b VDD VDD pfet
M16 n10 f n9 VDD pfet
M17 n7 g n10 VDD pfet
M18 n12 h n9 VDD pfet
M19 n7 i n12 VDD pfet
M20 n14 j n9 VDD pfet
M21 n7 k n14 VDD pfet
M22 n7 a VDD VDD pfet
A equação é :(a*(b*(c+d*(e+f))+g*h*i))
M1 n1 e GND GND nfet
M2 n1 f GND GND nfet
M3 n2 d n1 GND nfet
M4 n2 c GND GND nfet
M5 n7 b n2 GND nfet
M6 n4 g GND GND nfet
M7 n5 h n4 GND nfet
M8 n7 i n5 GND nfet
M9 n7 a n7 GND nfet
M10 n8 e VDD VDD pfet
M11 n9 f n8 VDD pfet
M12 n9 d VDD VDD pfet
M13 n10 c n9 VDD pfet
M14 n10 b VDD VDD pfet
M15 n7 g n10 VDD pfet
M16 n7 h n10 VDD pfet
M17 n7 i n10 VDD pfet
M18 n7 a VDD VDD pfet
